`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    02:31:07 02/11/2019 
// Design Name: 
// Module Name:    alu 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module alu (a,b,aluc,r,z); // 32-bit alu with a zero flag
input [31:0] a, b; // inputs: a, b
input [3:0] aluc;
output [31:0] r; // output: alu result // x 0 0 0 ADD
output z; // output: zero flag // x 1 0 0 SUB
wire [31:0] d_and = a & b; // x 0 0 1 AND
wire [31:0] d_or = a | b; // x 1 0 1 OR
wire [31:0] d_xor = a ^ b; // x 0 1 0 XOR
wire [31:0] d_lui = {b[15:0],16'h0}; // x 1 1 0 LUI
wire [31:0] d_and_or = aluc[2]? d_or : d_and; // 0 0 1 1 SLL
wire [31:0] d_xor_lui = aluc[2]? d_lui : d_xor; // 0 1 1 1 SRL
wire [31:0] d_as, d_sh; // 1 1 1 1 SRA
// addsub32 (a,b,sub, s);
addsub32 as32 (a,b,aluc[2],d_as); // add/sub
// shift (d,sa, right, arith, sh);
shift shifter (b,a[4:0],aluc[2],aluc[3],d_sh); // shift
// mux4x32 (a0, a1, a2, a3, s, y);
mux4x32 res (d_as,d_and_or,d_xor_lui,d_sh,aluc[1:0],r); // alu result
assign z = ~|r; // z = (r == 0)
endmodule